module contador_3bits(Clear, Clock, Tstep, Run, Resetn);

  /*
  Usado pela unidade de controle para saber em que etapa da instrução está.
   
  Ao receber Clear, volta para T0.
   
  Caso contrário, incrementa em cada borda de subida do clock.
  */

  input Clear, Clock, Run, Resetn;
  output reg [2:0] Tstep;
  reg Espera1ciclo_d = 0; // armazena o valor anterior de Espera1ciclo
  reg Resetn_d = 1;                   // armazena o valor anterior de Resetn
  reg Run_d = 0;                   // armazena o valor anterior de Run
  always @(posedge Clock)
    if (Clear && !Resetn) // se Clear for alto e Resetn for baixo, volta para T0
      begin
        Tstep <= 2'b0;
        Espera1ciclo_d <= 0; // atualiza Espera1ciclo_d para o próximo ciclo
      end
  /* else if (Run && !Run_d) // se Run for alto e Run_d for baixo, incrementa
    begin
      Tstep <= 2'b0;
      Run_d <= Run; // atualiza Run_d para o próximo ciclo
    end */
    /* else if (Espera1ciclo && !Espera1ciclo_d) // se Espera1ciclo for alto e Espera1ciclo_d for baixo, mantém Tstep
      begin
        Tstep <= Tstep;
        Espera1ciclo_d <= 1; // atualiza Espera1ciclo_d para o próximo ciclo
        $display("[%0t] linha 20 contador2bit Esperando um ciclo",$time);
      end */
    
    else if(Run)
      begin
        Tstep <= Tstep + 1'b1;
        Espera1ciclo_d <= 0; // atualiza Espera1ciclo_d para o próximo ciclo
      end
    else if (Resetn)
      begin
        // $display("[%0t] linha 20 contador2bit",$time);
        Tstep <= 2'b0; // Avaliar se coloca 11
      end
endmodule
module decode3_8bits(W, En, Y);

/*
   3bits to 8 bits decoder
   Transforma o campo XXX ou YYY
   da instrução em um sinal que pode ativar diretamente 
   um registrador específico (R0in, R1out, etc.). 
*/

  input [2:0] W;    // Codigo do registrador (campo XXX ou YYY da instrução)
  input En;         // Habilita o decodificador
  output [7:0] Y;  // Sinal de habilitação do registrador (R0in, R1out, etc.)
  reg [7:0] Y;
  always @(W or En)
    begin
      if (En == 1)
        case (W)
          3'b000:
            Y = 8'b1000_0000;
          3'b001:
            Y = 8'b0100_0000;
          3'b010:
            Y = 8'b0010_0000;
          3'b011:
            Y = 8'b0001_0000;
          3'b100:
            Y = 8'b0000_1000;
          3'b101:
            Y = 8'b0000_0100;
          3'b110:
            Y = 8'b0000_0010;
          3'b111:
            Y = 8'b0000_0001;
        endcase
      else
        Y = 8'b00000000;
    end
endmodule
// megafunction wizard: %RAM: 1-PORT%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altsyncram 

// ============================================================
// File Name: memoram.v
// Megafunction Name(s):
// 			altsyncram
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 13.0.1 Build 232 06/12/2013 SP 1 SJ Web Edition
// ************************************************************


//Copyright (C) 1991-2013 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
// synopsys translate_on
module memoram_dados (
	address,
	clock,
	data,
	wren,
	q);

	input	[5:0]  address;
	input	  clock;
	input	[15:0]  data;
	input	  wren;
	output	[15:0]  q;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri1	  clock;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire [15:0] sub_wire0;
	wire [15:0] q = sub_wire0[15:0];

	altsyncram	altsyncram_component (
				.address_a (address),
				.clock0 (clock),
				.data_a (data),
				.wren_a (wren),
				.q_a (sub_wire0),
				.aclr0 (1'b0),
				.aclr1 (1'b0),
				.address_b (1'b1),
				.addressstall_a (1'b0),
				.addressstall_b (1'b0),
				.byteena_a (1'b1),
				.byteena_b (1'b1),
				.clock1 (1'b1),
				.clocken0 (1'b1),
				.clocken1 (1'b1),
				.clocken2 (1'b1),
				.clocken3 (1'b1),
				.data_b (1'b1),
				.eccstatus (),
				.q_b (),
				.rden_a (1'b1),
				.rden_b (1'b1),
				.wren_b (1'b0));
	defparam
		altsyncram_component.clock_enable_input_a = "BYPASS",
		altsyncram_component.clock_enable_output_a = "BYPASS",
		//altsyncram_component.init_file = "./pratica1_Giovanni_Thales/memoria_pratica1.mif",
		altsyncram_component.intended_device_family = "Cyclone II",
		altsyncram_component.lpm_hint = "ENABLE_RUNTIME_MOD=NO",
		altsyncram_component.lpm_type = "altsyncram",
		altsyncram_component.numwords_a = 64,
		altsyncram_component.operation_mode = "SINGLE_PORT",
		altsyncram_component.outdata_aclr_a = "NONE",
		altsyncram_component.outdata_reg_a = "CLOCK0",
		altsyncram_component.power_up_uninitialized = "FALSE",
		altsyncram_component.ram_block_type = "M4K",
		altsyncram_component.widthad_a = 6,
		altsyncram_component.width_a = 16,
		altsyncram_component.width_byteena_a = 1, 
		altsyncram_component.init_file = "dados_pratica2_1.mif";


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: ADDRESSSTALL_A NUMERIC "0"
// Retrieval info: PRIVATE: AclrAddr NUMERIC "0"
// Retrieval info: PRIVATE: AclrByte NUMERIC "0"
// Retrieval info: PRIVATE: AclrData NUMERIC "0"
// Retrieval info: PRIVATE: AclrOutput NUMERIC "0"
// Retrieval info: PRIVATE: BYTE_ENABLE NUMERIC "0"
// Retrieval info: PRIVATE: BYTE_SIZE NUMERIC "8"
// Retrieval info: PRIVATE: BlankMemory NUMERIC "0"
// Retrieval info: PRIVATE: CLOCK_ENABLE_INPUT_A NUMERIC "0"
// Retrieval info: PRIVATE: CLOCK_ENABLE_OUTPUT_A NUMERIC "0"
// Retrieval info: PRIVATE: Clken NUMERIC "0"
// Retrieval info: PRIVATE: DataBusSeparated NUMERIC "1"
// Retrieval info: PRIVATE: IMPLEMENT_IN_LES NUMERIC "0"
// Retrieval info: PRIVATE: INIT_FILE_LAYOUT STRING "PORT_A"
// Retrieval info: PRIVATE: INIT_TO_SIM_X NUMERIC "0"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
// Retrieval info: PRIVATE: JTAG_ENABLED NUMERIC "0"
// Retrieval info: PRIVATE: JTAG_ID STRING "NONE"
// Retrieval info: PRIVATE: MAXIMUM_DEPTH NUMERIC "0"
// Retrieval info: PRIVATE: MIFfilename STRING "./pratica1_Giovanni_Thales/memoria_pratica1.mif"
// Retrieval info: PRIVATE: NUMWORDS_A NUMERIC "64"
// Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "2"
// Retrieval info: PRIVATE: READ_DURING_WRITE_MODE_PORT_A NUMERIC "3"
// Retrieval info: PRIVATE: RegAddr NUMERIC "1"
// Retrieval info: PRIVATE: RegData NUMERIC "1"
// Retrieval info: PRIVATE: RegOutput NUMERIC "1"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: SingleClock NUMERIC "1"
// Retrieval info: PRIVATE: UseDQRAM NUMERIC "1"
// Retrieval info: PRIVATE: WRCONTROL_ACLR_A NUMERIC "0"
// Retrieval info: PRIVATE: WidthAddr NUMERIC "6"
// Retrieval info: PRIVATE: WidthData NUMERIC "16"
// Retrieval info: PRIVATE: rden NUMERIC "0"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: CLOCK_ENABLE_INPUT_A STRING "BYPASS"
// Retrieval info: CONSTANT: CLOCK_ENABLE_OUTPUT_A STRING "BYPASS"
// Retrieval info: CONSTANT: INIT_FILE STRING "./pratica1_Giovanni_Thales/memoria_pratica1.mif"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
// Retrieval info: CONSTANT: LPM_HINT STRING "ENABLE_RUNTIME_MOD=NO"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altsyncram"
// Retrieval info: CONSTANT: NUMWORDS_A NUMERIC "64"
// Retrieval info: CONSTANT: OPERATION_MODE STRING "SINGLE_PORT"
// Retrieval info: CONSTANT: OUTDATA_ACLR_A STRING "NONE"
// Retrieval info: CONSTANT: OUTDATA_REG_A STRING "CLOCK0"
// Retrieval info: CONSTANT: POWER_UP_UNINITIALIZED STRING "FALSE"
// Retrieval info: CONSTANT: RAM_BLOCK_TYPE STRING "M4K"
// Retrieval info: CONSTANT: WIDTHAD_A NUMERIC "6"
// Retrieval info: CONSTANT: WIDTH_A NUMERIC "16"
// Retrieval info: CONSTANT: WIDTH_BYTEENA_A NUMERIC "1"
// Retrieval info: USED_PORT: address 0 0 6 0 INPUT NODEFVAL "address[5..0]"
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT VCC "clock"
// Retrieval info: USED_PORT: data 0 0 16 0 INPUT NODEFVAL "data[15..0]"
// Retrieval info: USED_PORT: q 0 0 16 0 OUTPUT NODEFVAL "q[15..0]"
// Retrieval info: USED_PORT: wren 0 0 0 0 INPUT NODEFVAL "wren"
// Retrieval info: CONNECT: @address_a 0 0 6 0 address 0 0 6 0
// Retrieval info: CONNECT: @clock0 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: @data_a 0 0 16 0 data 0 0 16 0
// Retrieval info: CONNECT: @wren_a 0 0 0 0 wren 0 0 0 0
// Retrieval info: CONNECT: q 0 0 16 0 @q_a 0 0 16 0
// Retrieval info: GEN_FILE: TYPE_NORMAL memoram.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL memoram.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL memoram.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL memoram.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL memoram_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL memoram_bb.v TRUE
// Retrieval info: LIB_FILE: altera_mf
// megafunction wizard: %RAM: 1-PORT%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altsyncram 

// ============================================================
// File Name: memoram.v
// Megafunction Name(s):
// 			altsyncram
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 13.0.1 Build 232 06/12/2013 SP 1 SJ Web Edition
// ************************************************************


//Copyright (C) 1991-2013 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
// synopsys translate_on
module memoram (
	address,
	clock,
	data,
	wren,
	q);

	input	[5:0]  address;
	input	  clock;
	input	[15:0]  data;
	input	  wren;
	output	[15:0]  q;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri1	  clock;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire [15:0] sub_wire0;
	wire [15:0] q = sub_wire0[15:0];

	altsyncram	altsyncram_component (
				.address_a (address),
				.clock0 (clock),
				.data_a (data),
				.wren_a (wren),
				.q_a (sub_wire0),
				.aclr0 (1'b0),
				.aclr1 (1'b0),
				.address_b (1'b1),
				.addressstall_a (1'b0),
				.addressstall_b (1'b0),
				.byteena_a (1'b1),
				.byteena_b (1'b1),
				.clock1 (1'b1),
				.clocken0 (1'b1),
				.clocken1 (1'b1),
				.clocken2 (1'b1),
				.clocken3 (1'b1),
				.data_b (1'b1),
				.eccstatus (),
				.q_b (),
				.rden_a (1'b1),
				.rden_b (1'b1),
				.wren_b (1'b0));
	defparam
		altsyncram_component.clock_enable_input_a = "BYPASS",
		altsyncram_component.clock_enable_output_a = "BYPASS",
		//altsyncram_component.init_file = "./pratica1_Giovanni_Thales/memoria_pratica1.mif",
		altsyncram_component.intended_device_family = "Cyclone II",
		altsyncram_component.lpm_hint = "ENABLE_RUNTIME_MOD=NO",
		altsyncram_component.lpm_type = "altsyncram",
		altsyncram_component.numwords_a = 64,
		altsyncram_component.operation_mode = "SINGLE_PORT",
		altsyncram_component.outdata_aclr_a = "NONE",
		altsyncram_component.outdata_reg_a = "CLOCK0",
		altsyncram_component.power_up_uninitialized = "FALSE",
		altsyncram_component.ram_block_type = "M4K",
		altsyncram_component.widthad_a = 6,
		altsyncram_component.width_a = 16,
		altsyncram_component.width_byteena_a = 1, 
		altsyncram_component.init_file = "instrucoes_pratica2_1.mif";


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: ADDRESSSTALL_A NUMERIC "0"
// Retrieval info: PRIVATE: AclrAddr NUMERIC "0"
// Retrieval info: PRIVATE: AclrByte NUMERIC "0"
// Retrieval info: PRIVATE: AclrData NUMERIC "0"
// Retrieval info: PRIVATE: AclrOutput NUMERIC "0"
// Retrieval info: PRIVATE: BYTE_ENABLE NUMERIC "0"
// Retrieval info: PRIVATE: BYTE_SIZE NUMERIC "8"
// Retrieval info: PRIVATE: BlankMemory NUMERIC "0"
// Retrieval info: PRIVATE: CLOCK_ENABLE_INPUT_A NUMERIC "0"
// Retrieval info: PRIVATE: CLOCK_ENABLE_OUTPUT_A NUMERIC "0"
// Retrieval info: PRIVATE: Clken NUMERIC "0"
// Retrieval info: PRIVATE: DataBusSeparated NUMERIC "1"
// Retrieval info: PRIVATE: IMPLEMENT_IN_LES NUMERIC "0"
// Retrieval info: PRIVATE: INIT_FILE_LAYOUT STRING "PORT_A"
// Retrieval info: PRIVATE: INIT_TO_SIM_X NUMERIC "0"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
// Retrieval info: PRIVATE: JTAG_ENABLED NUMERIC "0"
// Retrieval info: PRIVATE: JTAG_ID STRING "NONE"
// Retrieval info: PRIVATE: MAXIMUM_DEPTH NUMERIC "0"
// Retrieval info: PRIVATE: MIFfilename STRING "./pratica1_Giovanni_Thales/memoria_pratica1.mif"
// Retrieval info: PRIVATE: NUMWORDS_A NUMERIC "64"
// Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "2"
// Retrieval info: PRIVATE: READ_DURING_WRITE_MODE_PORT_A NUMERIC "3"
// Retrieval info: PRIVATE: RegAddr NUMERIC "1"
// Retrieval info: PRIVATE: RegData NUMERIC "1"
// Retrieval info: PRIVATE: RegOutput NUMERIC "1"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: SingleClock NUMERIC "1"
// Retrieval info: PRIVATE: UseDQRAM NUMERIC "1"
// Retrieval info: PRIVATE: WRCONTROL_ACLR_A NUMERIC "0"
// Retrieval info: PRIVATE: WidthAddr NUMERIC "6"
// Retrieval info: PRIVATE: WidthData NUMERIC "16"
// Retrieval info: PRIVATE: rden NUMERIC "0"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: CLOCK_ENABLE_INPUT_A STRING "BYPASS"
// Retrieval info: CONSTANT: CLOCK_ENABLE_OUTPUT_A STRING "BYPASS"
// Retrieval info: CONSTANT: INIT_FILE STRING "./pratica1_Giovanni_Thales/memoria_pratica1.mif"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
// Retrieval info: CONSTANT: LPM_HINT STRING "ENABLE_RUNTIME_MOD=NO"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altsyncram"
// Retrieval info: CONSTANT: NUMWORDS_A NUMERIC "64"
// Retrieval info: CONSTANT: OPERATION_MODE STRING "SINGLE_PORT"
// Retrieval info: CONSTANT: OUTDATA_ACLR_A STRING "NONE"
// Retrieval info: CONSTANT: OUTDATA_REG_A STRING "CLOCK0"
// Retrieval info: CONSTANT: POWER_UP_UNINITIALIZED STRING "FALSE"
// Retrieval info: CONSTANT: RAM_BLOCK_TYPE STRING "M4K"
// Retrieval info: CONSTANT: WIDTHAD_A NUMERIC "6"
// Retrieval info: CONSTANT: WIDTH_A NUMERIC "16"
// Retrieval info: CONSTANT: WIDTH_BYTEENA_A NUMERIC "1"
// Retrieval info: USED_PORT: address 0 0 6 0 INPUT NODEFVAL "address[5..0]"
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT VCC "clock"
// Retrieval info: USED_PORT: data 0 0 16 0 INPUT NODEFVAL "data[15..0]"
// Retrieval info: USED_PORT: q 0 0 16 0 OUTPUT NODEFVAL "q[15..0]"
// Retrieval info: USED_PORT: wren 0 0 0 0 INPUT NODEFVAL "wren"
// Retrieval info: CONNECT: @address_a 0 0 6 0 address 0 0 6 0
// Retrieval info: CONNECT: @clock0 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: @data_a 0 0 16 0 data 0 0 16 0
// Retrieval info: CONNECT: @wren_a 0 0 0 0 wren 0 0 0 0
// Retrieval info: CONNECT: q 0 0 16 0 @q_a 0 0 16 0
// Retrieval info: GEN_FILE: TYPE_NORMAL memoram.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL memoram.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL memoram.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL memoram.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL memoram_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL memoram_bb.v TRUE
// Retrieval info: LIB_FILE: altera_mf
module mux(
    input  wire [7:0]  Rout,          // seleção do registrador
    input  wire        Gout,          // habilita leitura de G
    input  wire        DINout,        // habilita leitura de DIN
    input  wire [15:0] R0out,
    input  wire [15:0] R1out,
    input  wire [15:0] R2out,
    input  wire [15:0] R3out,
    input  wire [15:0] R4out,
    input  wire [15:0] R5out,
    input  wire [15:0] R6out,
    input  wire [15:0] R7out,
    input  wire [15:0] Gout_data,
    input  wire [15:0] DINout_data,
    input  wire [15:0] Memout_data,  // dado de saída da memória
    input  wire        Memout,       // habilita leitura de Memout
    input  wire        Resetn,              // sinal de reset
    output reg  [15:0] BusWires
  );

  always @(DINout or Gout or Rout or Resetn or Memout)
    begin
      // Prioridade: DINout > Gout > Rout
      if (DINout)
        begin
          BusWires = DINout_data;
        end
      else if (Gout)
        begin
          BusWires = Gout_data;
        end
      else if (Resetn)
        begin
          BusWires = 16'b0;  // valor de reset no bus
        end
      else if (Memout)
        begin
          BusWires = Memout_data;  // dado de saída da memória
        end
      else
        begin
          case (Rout)
            8'b1000_0000:
              BusWires = R0out;
            8'b0100_0000:
              BusWires = R1out;
            8'b0010_0000:
              BusWires = R2out;
            8'b0001_0000:
              BusWires = R3out;
            8'b0000_1000:
              BusWires = R4out;
            8'b0000_0100:
              BusWires = R5out;
            8'b0000_0010:
              BusWires = R6out;
            8'b0000_0001:
              BusWires = R7out;
            default:
              BusWires = 16'bx;  // valor indefinido se nada selecionado
          endcase
        end
    end

endmodule
module processador_multiciclo (Resetn,
                                 Clock, Run, Done, BusWires, Rx_data, Ry_data, Tstep);

  /*
    
    Um processador multiciclo simples, com 8 registradores de 16 bits (R0 a R7), um registrador de 16 bits A, 
  um registrador de 16 bits G e uma ALU de soma/subtracao.
   
  Possui:
      -Um contador (Tstep) controla os ciclos de execucao (T1, T2, T3).
      -Um registrador de instrcao (IR) guarda a instruo atual.
      -Sinais de controle s£o gerados dependendo da etapa (Tstep_Q) e do opcode (I).
      -Registradores (R0 a R7, A, G) e a ALU (soma/subtrao) s£o instanciados.
      -Um multiplexador define o valor presente no BusWires a cada momento.
      -Um case aninhado © usado para acionar os sinais corretos de controle a cada T1/T2/T3.
  */

  /*
  killmodelsim;vlog processador_multiciclo.v registrador.v registrador_IR.v mux.v unidade_controle.v contador_2bits.v;vsim -L altera work.processador_multiciclo
  */


  // input [15:0] DIN; // deve ser 000 000 001 para comecar
  input Resetn, Clock, Run;
  output Done;
  output wire [15:0] BusWires;
  // output reg [15:0] BusWires;


  // Variaveis para controle
  wire [9:0] Instrucao;
  output wire [2:0] Tstep; // 00=T0,01=T1,10=T2,11=T3
  wire W_D;
  wire Clear;
  wire IncrPc;

  // Para o mux
  wire [15:0] DIN;            // barramento de entrada de dados
  wire [7:0]  Rout, Rin;      // campo de seleo para os registradores
  wire [9:0]  IRout;          // Saida do registrador IR
  wire [15:0] R0out, R1out, R2out, R3out, R4out, R5out, R6out, R7out; // saida do registrador R0, R1, ..., R7
  wire [15:0] ARout;          // saida do registrador GOUT
  wire [15:0] GRout;          // saida do registrador GOUT
  wire [15:0] ADDRout;        // saida do registrador ADDR
  wire [15:0] Memout_data;        // saida do registrador ADDR
  wire [15:0] DOUTout;        // saida do registrador DOUT
  wire [15:0] Ulaout;         // saida da ULA
  wire [2:0]  Ulaop;           // operacao da Ula
  wire        IRin, Ain, Gin, ADDRin, DOUTin; // habilita escrita no IR, A, G, ADDR e DOUT
  wire        Gout;           // habilita leitura do registrador G
  wire        DINout;         // habilita a saida do barramento DIN
  wire        Memout;         // habilita a saida do barramento Memout  
  wire [15:0] BusWires_data;  // dados do barramento BusWires
  wire [5:0]  endereco_mem; // endereco da memoria de dados

  assign endereco_mem = ADDRout[5:0];
  assign Instrucao = IRout;

  // Variaveis inuteis
  wire [8:0] UnusedQ9;
  wire [15:0] UnusedQ16;
  wire [15:0] NumeroInstrucoesExecutadas;
  wire [3:0]  Opcode;

  assign Opcode = Instrucao[9:6]; // opcode III

  // Variaveis da simulacao FPGA
  wire [2:0] Rx = IRout[5:3];
  wire [2:0] Ry = IRout[2:0];
  output [15:0] Rx_data; // Dados do registrador Rx
  output [15:0] Ry_data; // Dados do registrador Ry
  reg [15:0] Rx_data_reg, Ry_data_reg;
  reg [15:0] LazyBusWires;
  reg [7:0] LazyRin;
  assign Rx_data = Rx_data_reg;
  assign Ry_data = Ry_data_reg;
  // assign BusWires = LazyBusWires;
  // assign Rin = LazyRin;


  // wire [8:0] useless_IR_out =

  memoram_dados Memoria_Dados (
            .address(endereco_mem), // tem 64 enderecos,
            // .address(6'b001010), // tem 64 enderecos,
            .clock(Clock),
            .data(DOUTout),
            .wren(W_D),
            .q(Memout_data)
          );

  memoram Memoria_instrucao (
            .address(R7out[5:0]), // tem 64 enderecos,
            // .address(6'b000_000), // tem 64 enderecos,
            .clock(Clock),
            .data(DOUTout),
            .wren(1'b0), // nao escreve na memoria de instrucao nunca
            .q(DIN)
          );

  registrador_IR IR (
                   .R     (DIN[9:0]),          // entrada de dados (dado a ser escrito)
                   .Rin   (IRin),              // habilita escrita no registrador
                   .Clock (Clock),             // sinal de clock
                   .Resetn(Resetn),         // sinal de reset
                   .Q     (IRout)              // saida Inutil
                 );

  registrador_PC R7(
				.R      (BusWires     ),
				.Rin    (Rin[0]       ),
				.Clock  (Clock        ),
				.Resetn (Resetn       ),
				.IncrPc (IncrPc       ),
				.Q      (R7out        )
			 );

  registrador ADDR (
                .R    (BusWires),         // entrada de dados (dado a ser escrito)
                .Rin  (ADDRin),           // habilita escrita no registrador
                .Resetn(Resetn),        // sinal de reset
                .Clock(Clock),            // sinal de clock
                .Q    (ADDRout)           // saida Inutil
              );

  registrador DOUT (
                .R    (BusWires),         // entrada de dados (dado a ser escrito)
                .Rin  (DOUTin),            // habilita escrita no registrador
                .Resetn(Resetn),          // sinal de reset
                .Clock(Clock),             // sinal de clock
                .Q    (DOUTout)          // saida Inutil
              );

 /*  contaInstrucao u_contaInstrucao(
      .Resetn (Resetn ),
      .Done   (Done   ),
      .Q      (NumeroInstrucoesExecutadas      )
  ); */
  
  registrador R0 (
                .R    (BusWires),   // entrada de dados
                .Rin  (Rin[7]),    // habilita escrita
                .Clock(Clock),       // sinal de clock
                .Resetn(Resetn),     // sinal de reset
                .Q    (R0out)   // saida registrada
              );

  registrador R1 (
                .R    (BusWires),   // entrada de dados
                .Rin  (Rin[6]),    // habilita escrita
                .Clock(Clock),       // sinal de clock
                .Resetn(Resetn),     // sinal de reset
                .Q    (R1out)   // saida registrada
              );

  registrador R2 (
                .R    (BusWires),   // entrada de dados
                .Rin  (Rin[5]),    // habilita escrita
                .Clock(Clock),       // sinal de clock
                .Resetn(Resetn),     // sinal de reset
                .Q    (R2out)   // saida registrada
              );

  registrador R3 (
                .R    (BusWires),   // entrada de dados
                .Rin  (Rin[4]),    // habilita escrita
                .Clock(Clock),       // sinal de clock
                .Resetn(Resetn),     // sinal de reset
                .Q    (R3out)   // saida registrada
              );

  registrador R4 (
                .R    (BusWires),   // entrada de dados
                .Rin  (Rin[3]),    // habilita escrita
                .Clock(Clock),       // sinal de clock
                .Resetn(Resetn),     // sinal de reset
                .Q    (R4out)   // saida registrada
              );

  registrador R5 (
                .R    (BusWires),   // entrada de dados
                .Rin  (Rin[2]),    // habilita escrita
                .Clock(Clock),       // sinal de clock
                .Resetn(Resetn),     // sinal de reset
                .Q    (R5out)   // saida registrada
              );

  // Registrador SP
  registrador_SP R6 (
                .R    (BusWires),   // entrada de dados
                .Rin  (Rin[1]),    // habilita escrita
                .Clock(Clock),       // sinal de clock
                .Resetn(Resetn),     // sinal de reset
                .Q    (R6out)   // saida registrada
              );

  registrador A (
                .R    (BusWires),   // entrada de dados
                .Rin  (Ain),        // habilita escrita
                .Clock(Clock),      // sinal de clock
                .Resetn(Resetn),     // sinal de reset
                .Q    (ARout)        // saida registrada
              );

  registrador G (
                .R    (Ulaout),   // entrada de dados
                .Rin  (Gin),       // habilita escrita
                .Clock(Clock),       // sinal de clock
                .Resetn(Resetn),     // sinal de reset
                .Q    (GRout)   // saida registrada
              );

  contador_3bits u_contador_3bits(
                   .Clear     (Clear ),
                   .Clock     (Clock ),
                   .Run       (Run   ),
                   .Resetn    (Resetn),
                   .Tstep     (Tstep)
                 );

  unidade_controle u_unidade_controle(
                     .Instrucao (Instrucao ),
                     .Tstep     (Tstep     ),
                     .IncrPc    (IncrPc    ),
                     .Clock     (Clock     ),
                     .W_D       (W_D       ),
                     .ADDRin    (ADDRin    ),
                     .DOUTin    (DOUTin    ),
                     .Run       (Run       ),
                     .Resetn    (Resetn    ),
                     .Clear     (Clear     ),
                     .GRout     (GRout     ),
                     .IRin      (IRin      ),
                     .Rin       (Rin       ),
                     .Rout      (Rout      ),
                     .Ain       (Ain       ),
                     .Gin       (Gin       ),
                     .Gout      (Gout      ),
                     .Ulaop     (Ulaop     ),
                     .DINout    (DINout    ),
                     .Memout    (Memout    ),        
                     .Done      (Done      )
                   );

  mux u_mux(
        .Rout        (Rout        ),
        .Resetn      (Resetn      ),
        .R0out       (R0out       ),
        .R1out       (R1out       ),
        .R2out       (R2out       ),
        .R3out       (R3out       ),
        .R4out       (R4out       ),
        .R5out       (R5out       ),
        .R6out       (R6out       ),
        .R7out       (R7out       ),
        .Gout        (Gout        ),  // Habilita colocar dados do registrador G no barramento BusWires
        .Gout_data   (GRout       ),  // Dados G para colocar no barramento BusWires DIN
        .DINout      (DINout      ),  // Habilita a saida do barramento DIN
        .DINout_data (DIN),           // Dados DIN para colocar no barramento BusWires DIN
        .Memout_data (Memout_data),   // Dados da Memoria de Dados para colocar no barramento BusWires
        .Memout      (Memout),        // Habilita a saida do barramento Memout
        .BusWires    (BusWires)
      );

  ula u_ula(
        .A        (ARout      ), // saida do registrador A
        .BusWires (BusWires   ),
        .Ulaop    (Ulaop      ),       // operao da ULA (soma ou subtrao)
        .Q        (Ulaout     ) // saida da ULA
      );

  assign Rx_data = Rx_data_reg;
  assign Ry_data = Ry_data_reg;

  always @(Clock)
    begin
      case (Rx)
        3'b000:
          Rx_data_reg = R0out;
        3'b001:
          Rx_data_reg = R1out;
        3'b010:
          Rx_data_reg = R2out;
        3'b011:
          Rx_data_reg = R3out;
        3'b100:
          Rx_data_reg = R4out;
        3'b101:
          Rx_data_reg = R5out;
        3'b110:
          Rx_data_reg = R6out;
        3'b111:
          Rx_data_reg = R7out;
      endcase

      case (Ry)
        3'b000:
          Ry_data_reg = R0out;
        3'b001:
          Ry_data_reg = R1out;
        3'b010:
          Ry_data_reg = R2out;
        3'b011:
          Ry_data_reg = R3out;
        3'b100:
          Ry_data_reg = R4out;
        3'b101:
          Ry_data_reg = R5out;
        3'b110:
          Ry_data_reg = R6out;
        3'b111:
          Ry_data_reg = R7out;
      endcase
    end




  /*
  killmodelsim;
  vlog processador_multiciclo.v registrador.v registrador_IR.v mux.v unidade_controle.v contador_2bits.v;
  vsim -L altera work.processador_multiciclo
  */


endmodule
module registrador_IR(R, Rin, Clock, Resetn, Q);
  // Modulo que representa um registrador de 16 bits que quando habilitado
  // armazena o valor Rin na entrada R. O valor armazenado é lido na

  // inputs
  input [9:0] R; // entrada de dados
  input Rin, Clock, Resetn; // Rin habilita escrita, Clock é o clock do processador, Resetn é o reset

  // outputs
  output reg [9:0] Q; // valor armazenado

  // reg [8:0] Q;
  always @(negedge Clock)
    begin
      if (Rin)
        begin
          // $display("[%0t] quero ve-la sorrir, Rin = %0d, R = %0d",$time, Rin, R);
          Q <= R; // armazena o valor de R no registrador Q
        end
      else if (Resetn)
        Q <= 9'd0; // Reseta o registrador Q para 0
    end

endmodule
module registrador_PC(R, IncrPc, Rin, Clock, Resetn, Q);
  // Modulo que representa um registrador de 16 bits que quando habilitado
  // armazena o valor Rin na entrada R. O valor armazenado é lido na

  // inputs
  input [15:0] R;
  input Rin, Clock, Resetn, IncrPc;

  // outputs
  output [15:0] Q; // valor armazenado

  reg [15:0] Q;
  // always @(negedge Clock or  Resetn or posedge IncrPc)
  always @(negedge Clock)
    begin
      if (Resetn)
        Q <= 16'd0;                         // Reset síncrono ativo em 1
      else if (Rin)
        Q <= R;                             // Load direto se Rin = 1
      else if (IncrPc)
        Q <= Q + 1;                         // Incrementa PC se habilitado
    end
endmodule
module registrador_SP(R, Rin, Clock, Resetn, Q);
  // Modulo que representa um registrador de 16 bits que quando habilitado
  // armazena o valor Rin na entrada R. O valor armazenado é lido na

  // inputs
  input [15:0] R;
  input Rin, Clock, Resetn;

  // outputs
  output [15:0] Q; // valor armazenado

  reg [15:0] Q;
  always @(negedge Clock)
    if (Rin && !Resetn) // se Rin for alto e Resetn for baixo, armazena R
      Q <= R;
    else if (Resetn)
      Q <= 16'd64; // Reseta o registrador Q para o tamanho maximo de memoria
endmodule
module registrador(R, Rin, Clock, Resetn, Q);
  // Modulo que representa um registrador de 16 bits que quando habilitado
  // armazena o valor Rin na entrada R. O valor armazenado é lido na

  // inputs
  input [15:0] R;
  input Rin, Clock, Resetn;

  // outputs
  output [15:0] Q; // valor armazenado

  reg [15:0] Q;
  always @(negedge Clock)
    if (Rin && !Resetn) // se Rin for alto e Resetn for baixo, armazena R
      Q <= R;
    else if (Resetn)
      Q <= 16'd0;
endmodule
/*
 Rodando no vscode
 vlib work
 vlib altera
 
 vlog -work altera /home/gi/altera/13.0sp1/modelsim_ase/altera/verilog/src/altera_mf.v
 
 vlog hierarquia_memoria.v memoram.v tb_hierarquia_memoria.v
 
 vsim -L altera tb_hierarquia_memoria
 */`timescale 1 ps / 1 ps

module tb_memoram;

  // Entradas
  reg [5:0] address;
  reg Clock;
  reg [15:0] data;
  reg wren;

  // Saída
  wire [15:0] q;

  // Instancia o módulo da memória
  memoram uut (
            .address(address),
            .clock(Clock),
            .data(data),
            .wren(wren),
            .q(q)
          );

  // Geração de Clock (10ns período)
  always #50 Clock = ~Clock;

  // Estímulos
  initial
    begin
      $display("Iniciando Testbench...");

      // Inicializações
      Clock = 0;
      address = 6'd1;
      data = 0;
      wren = 0;


      // Aguarda alguns ciclos
      @(posedge Clock);
      #1;

      @(posedge Clock);
      #1;
      $display("[%0t] Lendo endereco 1,demorou dois ciclos",$time);
      $display("[%0t] Endereco = %0d, Data = %0b",$time, address, q);
      
      wren = 1; // Habilita escrita
      data = 16'd42; // Valor a ser escrito
      @(posedge Clock);
      #1;
      $display("[%0t] Escrevendo no endereco 1 o valor 42",$time);
      $display("[%0t] Endereco = %0d, Data = %0d",$time, address, q);
      
      wren = 0; // Desabilita escrita
      @(posedge Clock);
      #1;
      $display("[%0t] Lendo endereco 1",$time);
      $display("[%0t] Endereco = %0d, Data = %0d",$time, address, q);

      address = 6'd2; // Muda o endereço para 2
      @(posedge Clock);
      #1;
      $display("[%0t] Lendo endereco 2",$time);
      $display("[%0t] Endereco = %0d, Data = %0d",$time, address, q);
      
      @(posedge Clock);
      #1;
      $display("[%0t] Lendo endereco 2",$time);
      $display("[%0t] Endereco = %0d, Data = %0d",$time, address, q);

      

      // Leitura da primeira posicao (endereço 0)
      $display("[%0t] Lendo endereco 0",$time);
      address = 6'd0;
      #100;
      $display("[%0t] Endereco = %0d, Data = %0b",$time, address, q);

      // Escrita no endereco 0
      $display("[%0t] Escrevendo no endereco 0 o valor 1",$time);
      address = 6'd0;
      data = 16'd1;
      wren = 1;
      #100;
      $display("[%0t] Endereco = %0d, Data = %0b",$time, address, q);

      // Leitura do endereco 0
      $display("[%0t] Lendo endereco 0",$time);
      address = 6'd0;
      wren = 0; // Desabilita escrita
      #100;
      $display("[%0t] Endereco = %0d, Data = %0b",$time, address, q);
      
      $stop;

      // Escreve valor 0xAAAA no endereço 5
      // address = 6'd5;
      // data = 16'hAAAA;
      // wren = 1;
      // #100;

      // // Escreve valor 0x1234 no endereço 10
      // address = 6'd10;
      // data = 16'h1234;
      // #100;

      // // Escreve valor 0xFFFF no endereço 20
      // address = 6'd20;
      // data = 16'hFFFF;
      // #100;

      // // Desabilita escrita
      // wren = 0;

      // // Lê dos mesmos endereços com atraso de Clock
      // #100;
      // address = 6'd5;
      // #10;
      // $display("Endereco 5 = %h (esperado: AAAA)", q);

      // address = 6'd10;
      // #10;
      // $display("Endereco 10 = %h (esperado: 1234)", q);

      // address = 6'd20;
      // #10;
      // $display("Endereco 20 = %h (esperado: FFFF)", q);

      // $display("Testbench finalizado.");
      // $stop;
    end

endmodule
`timescale 1ps/1ps

module tb_processador;

  reg [15:0] DIN;
  reg [2:0] Opcode;          // Opcode III
  reg [5:3] Rx;              // Rx (destino/target)
  reg [8:6] Ry;              // Ry (fonte/source)
  wire [8:0] Instrucao; // Instrução completa
  reg Clock, Resetn, Run;
  wire Done;
  wire [2:0] Tstep; // Sinal de Tstep
  wire [15:0] BusWires;
  wire [15:0] Rx_data, Ry_data; // Dados dos registradores Rx e Ry

  // Instancia o processador

  processador_multiciclo uut (
                           .Resetn   (Resetn   ),
                           .Clock    (Clock    ),
                           .Run      (Run      ),
                           .Done     (Done     ),
                           .BusWires (BusWires ),
                           .Tstep    (Tstep    ),
                           .Rx_data  (Rx_data  ),
                           .Ry_data  (Ry_data  )
                         );



  assign Instrucao = uut.Instrucao; // Instrução completa
  // Clock gerado a cada 50ps


  integer detalhado = 1;
  always #50 Clock = ~Clock;



  integer mostra_teste1 = 1;
  integer mostra_teste2 = 1;
  integer mostra_teste3 = 1;
  integer mostra_teste4 = 1;
  integer mostra_teste5 = 1;
  integer mostra_teste6 = 1;
  integer mostra_teste7 = 1;
  integer mostra_teste8 = 1;
  integer mostra_teste9 = 1;
  integer mostra_teste10 = 1;
  integer mostra_teste11 = 1;
  integer mostra_teste12 = 1;
  integer mostra_teste13 = 1;
  integer mostra_teste14 = 1;
  integer mostra_teste15 = 1;

  initial
    begin
      // Inicialização
      Clock = 0;
      Resetn = 1;
      Run = 0;
      DIN = 16'b0;
      // Reset do processador

      // ------------------------------
      // T0 - Resetn dos registradores e sinais
      // ------------------------------
      // @(posedge Clock);
      // #1;
      @(posedge Clock);
      #1;
      $display("[%0t] Teste Resetn (mux, registradores, e outros sinais)",$time);
      $display("[%0t] BusWires = %0d, DIN = %0d, Tstep = %0d",$time, BusWires, uut.DIN, uut.Tstep);
      $display("[%0t] R1 = %0d R2 = %0d, .. R6 = %0d R7 = %0b",$time, uut.R1.Q, uut.R2.Q, uut.R6.Q, uut.R7.Q);
      $display("[%0t] IncrPc=%0d W_D=%0d ADDRin=%0d DOUTin=%0d",
               $time, uut.IncrPc, uut.W_D, uut.ADDRin, uut.DOUTin);
      $display("[%0t] Run=%0d Resetn=%0d Clear=%0d GRout=%0d",
               $time, uut.Run, uut.Resetn, uut.Clear, uut.GRout);
      $display("[%0t] IRin=%0d Rin=%b Rout=%b Ain=%0d",
               $time, uut.IRin, uut.Rin, uut.Rout, uut.Ain);
      $display("[%0t] Gin=%0d Gout=%0d Ulaop=%b DINout=%h",
               $time, uut.Gin, uut.Gout, uut.Ulaop, uut.DINout);
      $display("[%0t] Done=%0d",
               $time, uut.Done);
      $display("[%0t] Teste 0 Finalizado",$time);
      $display("--------------------------------------------------");


      Run = 1; // Ativa o Run
      Resetn = 0; // Desativa o reset

      // -----------------------------
      // T1 - mvi R2 1
      // -----------------------------
      if (mostra_teste1)
        begin
          $display("[%0t] Teste 1 instrucao mvi R2 1, R2 com o valor inicial %0d, Tstep = %0d", $time, uut.R2.Q, uut.Tstep);
          @(posedge Clock);
          #351;
          $display("[%0t] Ciclo 5 NEG_EDGE", $time);
          $display("[%0t]           IR = %10b, R2 = %0d Tstep = %0d", $time, uut.IR.Q, uut.R2.Q, uut.Tstep);
          if (detalhado)
            $display("[%0t] ESPERADO: IR = 0001010000, R2 = 1 Tstep = 4",$time);
          $display("[%0t] Teste mvi R2 1 concluido.", $time);
          $display("--------------------------------------------------");
        end

      // -----------------------------
      // T2 - mvi R4 10
      // -----------------------------
      if (mostra_teste2)
        begin
          $display("[%0t] Teste 2 instrucao mvi R4 10, R4 com o valor inicial %0d, Tstep = %0d", $time, uut.R4.Q, uut.Tstep);
          @(posedge Clock);
          #451;
          $display("[%0t] Ciclo 5 NEG_EDGE", $time);
          $display("[%0t]           IR = %10b, R4 = %0d Tstep = %0d", $time, uut.IR.Q, uut.R4.Q, uut.Tstep);
          if (detalhado)
            $display("[%0t] ESPERADO: IR = 0001100000, R4 = 10 Tstep = 4",$time);
          $display("[%0t] Teste mvi R4 10 concluido.", $time);
          $display("--------------------------------------------------");
        end

      // -----------------------------
      // T3 - mvi R0 4
      // -----------------------------
      if (mostra_teste3)
        begin
          $display("[%0t] Teste 3 instrucao mvi R0 4, R4 com o valor inicial %0d, Tstep = %0d", $time, uut.R0.Q, uut.Tstep);
          @(posedge Clock);
          #451;
          $display("[%0t] Ciclo 5 NEG_EDGE", $time);
          $display("[%0t]           IR = %10b, R0 = %0d Tstep = %0d", $time, uut.IR.Q, uut.R0.Q, uut.Tstep);
          if (detalhado)
            $display("[%0t] ESPERADO: IR = 0001000000, R0 = 4 Tstep = 4",$time);
          $display("[%0t] Teste mvi R0 4 concluido.", $time);
          $display("--------------------------------------------------");
        end

      // -----------------------------
      // T4 - MV R5 R0
      // -----------------------------
      if (mostra_teste4)
        begin
          $display("[%0t] Teste 4 instrucao mv R5, R0 R5 inicial = %0d, R0 inicial = %0d, Tstep = %0d", $time, uut.R5.Q, uut.R0.Q, uut.Tstep);
          @(posedge Clock);
          #351;
          $display("[%0t] Ciclo 4 NEG_EDGE", $time);
          $display("[%0t]           IR = %10b, R0 = %0d, R5 = %0d Tstep = %0d", $time, uut.IR.Q, uut.R5.Q, uut.R0.Q, uut.Tstep);
          if (detalhado)
            $display("[%0t] ESPERADO: IR = 0000101000, R0 = 4  R5 = 4 Tstep = 3",$time);
          $display("[%0t] Teste mv R0 R5 1 concluido.", $time);
          $display("--------------------------------------------------");
        end

      // -----------------------------
      // T5 - mvnz R3 R2
      // -----------------------------
      if (mostra_teste5)
        begin
          $display("[%0t] Teste 5 instrucao mvnz R3, R3 inicial = %0d, R2 inicial = %0d, Tstep = %0d", $time, uut.R3.Q, uut.R2.Q, uut.Tstep);
          @(posedge Clock);
          #351;
          $display("[%0t] Ciclo 4 NEG_EDGE", $time);
          $display("[%0t]           IR = %10b, R3 = %0d, R2 = %0d Tstep = %0d", $time, uut.IR.Q, uut.R3.Q, uut.R2.Q, uut.Tstep);
          if (detalhado)
            $display("[%0t] ESPERADO: IR = 0010011010, R3 = 0  R2 = 1 Tstep = 3",$time);
          $display("[%0t] Teste mvnz R3 R2 concluido.", $time);
          $display("--------------------------------------------------");
        end

      // -----------------------------
      // T6- ADD R4, R2
      // -----------------------------
      if (mostra_teste6)
        begin
          $display("[%0t] Teste 6 instrucao add R4, R2, R4 inicial = %0d, R2 inicial = %0d, Tstep = %0d", $time, uut.R4.Q, uut.R2.Q, uut.Tstep);
          @(posedge Clock);
          #551;
          $display("[%0t] Ciclo 4 NEG_EDGE", $time);
          $display("[%0t]           IR = %10b, R4 = %0d, R2 = %0d Tstep = %0d", $time, uut.IR.Q, uut.R4.Q, uut.R2.Q, uut.Tstep);
          if (detalhado)
            $display("[%0t] ESPERADO: IR = 0100100010, R4 = 11  R2 = 1 Tstep = 5",$time);
          $display("[%0t] Teste add R4, R2 concluido.", $time);
          $display("--------------------------------------------------");
        end

      // -----------------------------
      // T7- SUB R4, R2
      // -----------------------------
      if (mostra_teste7)
        begin
          $display("[%0t] Teste 7 instrucao sub R4, R2, R4 inicial = %0d, R2 inicial = %0d, Tstep = %0d", $time, uut.R4.Q, uut.R2.Q, uut.Tstep);
          @(posedge Clock);
          #551;
          $display("[%0t] Ciclo 5 NEG_EDGE", $time);
          $display("[%0t]           IR = %10b, R4 = %0d, R2 = %0d Tstep = %0d", $time, uut.IR.Q, uut.R4.Q, uut.R2.Q, uut.Tstep);
          if (detalhado)
            $display("[%0t] ESPERADO: IR = 0100100010, R4 = 10  R2 = 1 Tstep = 5",$time);
          $display("[%0t] Teste sub R4, R2 concluido.", $time);
          $display("--------------------------------------------------");
        end

      // -----------------------------
      // T8 - SLT R1, R2
      // -----------------------------
      if (mostra_teste8)
        begin
          $display("[%0t] Teste 8 instrucao slt R1, R2, R1 inicial = %0d, R2 inicial = %0d, Tstep = %0d", $time, uut.R1.Q, uut.R2.Q, uut.Tstep);
          @(posedge Clock);
          #551;
          $display("[%0t] Ciclo 5 NEG_EDGE", $time);
          $display("[%0t]           IR = %10b, R1 = %0d, R2 = %0d Tstep = %0d", $time, uut.IR.Q, uut.R1.Q, uut.R2.Q, uut.Tstep);
          if (detalhado)
            $display("[%0t] ESPERADO: IR = 0100100010, R1 = 1  R2 = 4 Tstep = 5",$time);
          $display("[%0t] Teste slt R1, R2 concluido.", $time);
          $display("--------------------------------------------------");
        end

      // -----------------------------
      // T9 - LD R2, R1
      // -----------------------------
      if (mostra_teste9)
        begin
          $display("[%0t] Teste 9 instrucao LD R2, R1, R2 inicial = %0d, R1 inicial = %0d, Tstep = %0d", $time, uut.R2.Q, uut.R1.Q, uut.Tstep);
          @(posedge Clock);
          #551;
          $display("[%0t] Ciclo 5 NEG_EDGE", $time);
          $display("[%0t]           IR = %10b, R2 = %0d, R1 = %0d Tstep = %0d", $time, uut.IR.Q, uut.R2.Q, uut.R1.Q, uut.Tstep);
          if (detalhado)
            $display("[%0t] ESPERADO: IR = 0101001010, R2 = 2  R1 = 1 Tstep = 5",$time);
          $display("[%0t] Teste LD R2, R1 concluido.", $time);
          $display("--------------------------------------------------");
        end

      // ------------------------------
      // T10 - ST R1, R0 MODIFIQUEI CONTEUDO DE R1
      // ------------------------------
      if (mostra_teste10)
        begin
          uut.R1.Q = 16'd10; // R1 = 10
          $display("[%0t] Teste 10 instrucao ST R1, R0, R1 inicial = %0d, R0 inicial = %0d, Tstep = %0d", $time, uut.R1.Q, uut.R0.Q, uut.Tstep);
          @(posedge Clock);
          #451;
          $display("[%0t] Ciclo 5 NEG_EDGE", $time);
          $display("[%0t]           IR = %10b, R1 = %0d, R0 = %0d Tstep = %0d", $time, uut.IR.Q, uut.R1.Q, uut.R0.Q, uut.Tstep);
          if (detalhado)
            $display("[%0t] ESPERADO: IR = 0100100010, R1 = 10  R0 = 4 Tstep = 5",$time);
          $display("[%0t] Teste ST R1, R0 concluido.", $time);
          $display("--------------------------------------------------");
        end

      // ------------------------------
      // T11 - LD R3, R0
      // ------------------------------
      if (mostra_teste11)
        begin
          $display("[%0t] Teste 11 instrucao LD R3, R0, R3 inicial = %0d, R0 inicial = %0d, Tstep = %0d", $time, uut.R3.Q, uut.R0.Q, uut.Tstep);
          @(posedge Clock);
          #551;
          $display("[%0t] Ciclo 5 NEG_EDGE", $time);
          $display("[%0t]           IR = %10b, R3 = %0d, R0 = %0d Tstep = %0d", $time, uut.IR.Q, uut.R3.Q, uut.R0.Q, uut.Tstep);
          if (detalhado)
            $display("[%0t] ESPERADO: IR = 0101001010, R3 = 2  R0 = 1 Tstep = 5",$time);
          $display("[%0t] Teste LD R3, R0 concluido.", $time);
          $display("--------------------------------------------------");
        end

      // ------------------------------
      // T12 - PUSH R0
      // ------------------------------
      if (mostra_teste12)
        begin
          $display("[%0t] Teste 12 instrucao PUSH R0, R0 inicial = %0d, Tstep = %0d", $time, uut.R0.Q, uut.Tstep);
          @(posedge Clock);
          #551;
          $display("[%0t] Ciclo 5 NEG_EDGE", $time);
          $display("[%0t]           IR = %10b, R0 = %0d Tstep = %0d", $time, uut.IR.Q, uut.R0.Q, uut.Tstep);
          if (detalhado)
            $display("[%0t] ESPERADO: IR = 0101001010, R0 = 2 Tstep = 5",$time);
          $display("[%0t] Teste PUSH R0 concluido.", $time);
          $display("--------------------------------------------------");
        end

      // ------------------------------
      // T13 - LD R3, R6 - 4 MODIFIQUEI CONTEUDO DE R6
      // ------------------------------
      if (mostra_teste13)
        begin
          uut.R6.Q = 16'd60; // R2 = 2
          $display("[%0t] Teste 13 instrucao LD R3, R6, R3 inicial = %0d, R6 inicial = %0d, Tstep = %0d", $time, uut.R3.Q, uut.R6.Q, uut.Tstep);
          @(posedge Clock);
          #551;
          $display("[%0t] Ciclo 5 NEG_EDGE", $time);
          $display("[%0t]           IR = %10b, R3 = %0d, R6 = %0d Tstep = %0d", $time, uut.IR.Q, uut.R3.Q, uut.R6.Q, uut.Tstep);
          if (detalhado)
            $display("[%0t] ESPERADO: IR = 0101001010, R3 = 2  R6 = 1 Tstep = 5",$time);
          $display("[%0t] Teste LD R3, R6 concluido.", $time);
          $display("--------------------------------------------------");
        end

      // ------------------------------
      // T13 - POP R6 - 4 MODIFIQUEI CONTEUDO DE R6
      // ------------------------------
      if (mostra_teste14)
        begin
          uut.R6.Q = 16'd60; // R2 = 2
          $display("[%0t] Teste 14 instrucao POP R2, R2 inicial = %0d, Tstep = %0d", $time, uut.R2.Q, uut.Tstep);
          @(posedge Clock);
          #651;
          $display("[%0t] Ciclo 5 NEG_EDGE", $time);
          $display("[%0t]           IR = %10b, R2 = %0d Tstep = %0d", $time, uut.IR.Q, uut.R2.Q, uut.Tstep);
          if (detalhado)
            $display("[%0t] ESPERADO: IR = 0101001010, R2 = 2 Tstep = 5",$time);
          $display("[%0t] Teste POP R2 concluido.", $time);
          $display("--------------------------------------------------");
        end


      #300;
      $stop;

      // ------------------------------
      // T11 - ST R1, R0
      // ------------------------------

    end


  // Testes do AVA
  task teste_mvi_R2_1;
    begin
      Opcode = 3'b001; // mvi
      Rx = 3'b010;     // R2
      Ry = 3'b000;     // R0
      uut.R2.Q = 16'd0; // R0 = 11
      //uut.R1.Q = 16'd10; // R1 = 10
      DIN = {6'b000_000, Opcode, Rx, Ry}; // Formando a instrução: 000 001 010
    end
  endtask

  task teste_mvi_R4_10;
    begin
      Opcode = 3'b001; // mvi
      Rx = 3'b100;     // R0
      Ry = 3'b000;     // zzz
      uut.R4.Q = 16'd0; // R0 = 11
      //uut.R1.Q = 16'd10; // R1 = 10
      DIN = {6'b000_000, Opcode, Rx, Ry}; // Formando a instrução: 000 001 000
    end
  endtask

  task teste_mv_R5_R7;
    begin
      Opcode = 3'b000; // mvi
      Rx = 3'b101;     // R0
      Ry = 3'b111;     // zzz
      uut.R5.Q = 16'd1; // R0 = 11
      uut.R7.Q = 16'd2; // R0 = 11
      //uut.R1.Q = 16'd10; // R1 = 10
      DIN = {6'b000_000, Opcode, Rx, Ry}; // Formando a instrução: 000 001 000
    end
  endtask

  task teste_sub_R4_R2;
    begin
      Opcode = 3'b011; // sub
      Rx = 3'b100;     // R4
      Ry = 3'b010;     // R2
      uut.R4.Q = 16'd10; // R4 = 10
      uut.R2.Q = 16'd6; // R2 = 6
      DIN = {6'b000_000, Opcode, Rx, Ry}; // Formando a instrução: 000 001 000
    end
  endtask

  task teste_mvnz_R7_R5;
    begin
      Opcode = 3'b100; // mvnz
      Rx = 3'b111;     // R7
      Ry = 3'b101;     // R5
      uut.R7.Q = 16'd0; // R7 = 0
      uut.R5.Q = 16'd0; // R5 = 0
      uut.G.Q  = 16'd4; // G = 4
      DIN = {6'b000_000, Opcode, Rx, Ry}; // Formando a instrução: 000 001 000
    end
  endtask


  // Testes Internos

  task teste_mv_R0_R1;
    begin
      Opcode = 3'b000; // mv
      Rx = 3'b000;     // R0
      Ry = 3'b001;     // R1
      uut.R0.Q = 16'd11; // R0 = 11
      uut.R1.Q = 16'd10; // R1 = 10
      DIN = {6'b000_000, Opcode, Rx, Ry}; // Formando a instrução: 000 001 000
    end
  endtask

  task teste_mvi_R0_5;
    begin
      Opcode = 3'b001; // mv
      Rx = 3'b000;     // R0
      Ry = 3'b001;     // R1
      uut.R0.Q = 16'd11; // R0 = 11
      uut.R1.Q = 16'd10; // R1 = 10
      DIN = {6'b000_000, Opcode, Rx, Ry}; // Formando a instrução: 000 001 000
    end
  endtask

  task teste_sub_R1_R0;
    begin
      Opcode = 3'b011; // sub
      Rx = 3'b001;     // R1
      Ry = 3'b000;     // R0
      uut.R0.Q = 16'd5; // R0 = 11
      uut.R1.Q = 16'd10; // R1 = 10
      DIN = {6'b000_000, Opcode, Rx, Ry}; // Formando a instrução: 000 001 000
    end
  endtask

  task teste1_mvnz_R0_R1;
    begin
      Opcode = 3'b100; // mvnz
      Rx = 3'b000;     // R0
      Ry = 3'b001;     // R1
      uut.R0.Q = 16'd11; // R0 = 11
      uut.R1.Q = 16'd10; // R1 = 10
      uut.G.Q  = 16'd0;  // G = 0
      DIN = {6'b000_000, Opcode, Rx, Ry}; // Formando a instrução: 000 001 000
    end
  endtask

  task teste2_mvnz_R0_R1;
    begin
      Opcode = 3'b100; // mvnz
      Rx = 3'b000;     // R0
      Ry = 3'b001;     // R1
      uut.R0.Q = 16'd11; // R0 = 11
      uut.R1.Q = 16'd10; // R1 = 10
      uut.G.Q  = 16'd5;  // G = 0
      DIN = {6'b000_000, Opcode, Rx, Ry}; // Formando a instrução: 000 001 000
    end
  endtask



  task cabecalho_teste(input integer numero_task);
    begin
      $display("--------------------------------------------------");
      $display("[%0t] Teste %0d", $time, numero_task);
      $display("--------------------------------------------------");
    end
  endtask

  integer disp_sinais = 1;
  task meio_teste_1_ciclo;
    begin
      if (disp_sinais)
        $display("[%0t] Clock: %b, Resetn: %b, Run: %b, DIN: %b",$time, Clock, Resetn, Run, DIN);
      $display("[%0t] Barramento: %b, Tempo_Instrucao = %0d",$time, BusWires, uut.Tstep);
      $display("[%0t] Done: %b",$time, Done);
    end
  endtask

  /*
    always @(posedge Clock)
      begin
        counter_clock_cycle = counter_clock_cycle + 1;
        // $display("[%0t] Counter_Clock_Cycle ",$time);
        case (counter_clock_cycle)
          1:
            begin
              // Opcode = 3'b001; // mvi R0 5
              // Rx = 3'b000;     // R0
              // Ry = 3'b001;     // R1
              // uut.R0.Q = 16'd11; // R0 = 11
              // uut.R1.Q = 16'd10; // R1 = 10
              // DIN = {6'b000_000, Opcode, Rx, Ry}; // Formando a instrução: 000 001 000
              // cabecalho_teste(2);
              // Run = 1; // Agendado ja no inicio do ciclo
              // $display("[%0t] instrucao = %3b_%3b_%3b = mv R0 R1 000_000_001", $time, Instrucao[8:6], Instrucao[5:3], Instrucao[2:0]);
            end
   
   
        endcase
   
      end
  */


endmodule





/*
1 Ciclo em verilog
1. Avaliacao de condicoes, always, if,  e sinais agendados ( PROIBIDO USAR, ex: #2, se nao nao funciona FPGA)...
2. Blocking e Non Blocking, (SO use BLOCKING em logica dentro dos blocos),
3. Atribuicao dos Non Blocking Variaveis externas, sempre usar Non Blocking
 
clear;vsim -c -do vlog_terminal_tb_proc.do
killmodelsim;vsim -do vlog_wave_tb_proc.do 
alias killmodelsim='ps aux | grep '\''intelFPGA/20.1/'\'' | grep -v grep | awk '\''{print $2}'\'' | xargs kill -9'
*/
module ula(A, BusWires, Ulaop, Q);
  input [15:0] A, BusWires;
  input [2:0] Ulaop; // 2 bits para selecionar a operação da ULA
  output reg [15:0] Q; // Saída da ULA
  always @(A or BusWires or Ulaop)
    begin
      case (Ulaop)
        3'b000: // Adição
          Q <= A + BusWires;
        3'b001: // Subtração
          Q <= A - BusWires;
        3'b010: // SLT
          Q <= (A < BusWires) ? 16'd1 : 16'd0; // Set Less Than
        3'b011: // CMP
          Q <= (A == BusWires) ? 16'd1 : 16'd0; // Compare
        3'b100: // Soma 4
          Q <= BusWires + 16'd4; // Adição de 4
        3'b101: // Subtrai 4
          Q <= BusWires - 16'd4; // Subtração de 4
      endcase
    end
endmodule
// grupo 4
module unidade_controle (
    Instrucao,       // opcode III
    Tstep,   // 00=T0,01=T1,10=T2,11=T3
    Run,     // start instruction
    Clear,   // limpa contador de Tstep
    IncrPc, // incrementa PC
    GRout,   // saída do registrador G
    Memout,  // saída da memória
    IRin,    // carrega IR
    Rin,     // habilita escrita em R0..R7
    Rout,    // habilita leitura de R0..R7
    ADDRin, // habilita escrita no barramento
    DOUTin, // habilita escrita no barramento
    Ain,     // carrega registrador A
    Gin,     // carrega registrador G
    Gout,    // lê registrador G
    W_D, // habilita escrita no barramento
    Resetn,  // recomecar da primeira instrucao
    Ulaop,  // escolhe subtração na ALU
    DINout,  // coloca DIN no barramento
    Clock,
    Done     // instrucao concluída
  );

  parameter mv   = 4'b0000; // mv Rx,Ry
  parameter mvi  = 4'b0001; // mvi Rx,imediato
  parameter mvnz = 4'b0010; // mvnz Rx,Ry

  parameter add  = 4'b0011; // add Rx,Ry
  parameter sub  = 4'b0100; // sub Rx,Ry
  parameter slt  = 4'b0101; // slt Rx,Ry
  parameter cmp  = 4'b0110; // cmp Rx,Ry

  parameter ld   = 4'b0111; // ld Rx,imediato
  parameter st   = 4'b1000; // st Rx,imediato
  parameter push = 4'b1001; // push Rx
  parameter pop  = 4'b1010; // pop Rx

  /*
   contador_2bits u_contador_2bits(
    .Clear (Clear ),
    .Clock (Clock ),
    .Q     (Tstep )
  );
  */

  // inputs
  input  wire       Clock;      // clock do processador
  input  wire [9:0] Instrucao;  // opcode III CONECTA com o memoram
  input  wire [2:0] Tstep;      // 00=T0,01=T1,10=T2,11=T3
  input  wire       Run;        // start instruction
  input  wire       Resetn;     // recomecar da primeira instrucao
  input  wire [15:0] GRout;       // saída do registrador G

  // outputs
  output reg        IncrPc;
  output reg        W_D;
  output reg        Clear;   // limpa contador de Tstep
  output reg        IRin;    // carrega IR
  output reg        ADDRin;                // habilita escrita no barramento
  output reg        DOUTin;                // habilita escrita no barramento
  // output wire [7:0]  Rin;     // habilita escrita em R0..R7
  // output wire [7:0]  Rout;    // habilita leitura de R0..R7
  output reg [7:0]  Rin;     // habilita escrita em R0..R7
  output reg [7:0]  Rout;    // habilita leitura de R0..R7
  output reg        Ain;     // carrega registrador A
  output reg        Gin;     // carrega registrador G
  output reg        Gout;    // lê registrador G
  output reg        Memout;   // le da memoria
  output reg [2:0]  Ulaop;  // escolhe subtração ou adicao na ALU
  output reg        DINout;  // coloca DIN no barramento
  output reg        Done;    // instrucao concluída

  // Variaveis
  reg Run_d = 0;                   // armazena o valor anterior de Run
  reg Resetn_d = 1;                   // armazena o valor anterior de Run
  reg En;                     // habilita o decodificador
  wire [3:0] opcode;           // opcode III
  wire [5:3] Rx;              // campo destino
  wire [8:6] Ry;              // campo fonte
  wire [7:0] Wire_Rin;        // campo de seleção para os registradores
  wire [7:0] Wire_Rout;       // campo de seleção para os registradores


  // Instanciacoes
  assign Ry     = Instrucao[2:0]; // campo fonte   (quem fornece o dado)
  assign Rx     = Instrucao[5:3]; // campo destino (quem fica com o dado fornecido)
  assign opcode = Instrucao[9:6]; // opcode IIII
  //Run_d = 0; // inicializa Run_d



  decode3_8bits Rx_decode3_8bits(
                  .W  (Rx  ), // campo XXX ou YYY da instrução
                  .En (1'b1 ), // Habilita o decodificador
                  .Y  (Wire_Rin ) // Sinal de habilitação do registrador (R0in, R1out, etc.)
                );
  // Logica do registrador destino (out)
  decode3_8bits Ry_decode3_8bits(
                  .W  (Ry  ),
                  .En (1'b1 ), // Habilita o decodificador
                  .Y  (Wire_Rout ) // Sinal de habilitação do registrador (R0in, R1out, etc.)
                );

  // always @(Tstep or Run or Resetn) // or Resetn
  always @(Tstep or Resetn) // or Resetn
    begin
      /* Todos os sinais mudados aqui, devem ser alterados com <=, pq se nao fica com 0 pq eh non blocking*/
      if (Resetn && !Run ) // Reset ativo em nível baixo
        begin
          Resetn_d <= 1; // reseta o valor de Resetn_d
          Run_d   <= 0; // reseta Run_d
          Clear   <= 1; // limpa o contador de Tstep
          IncrPc  <= 0; // não incrementa o PC
          W_D     <= 0; // não habilita escrita no barramento
          Clear   <= 1; // limpa o contador de Tstep
          IRin    <= 0; // não carrega IR
          Rin     <= 8'b0; // não habilita escrita em R0..R7
          Rout    <= 8'b0; // não habilita leitura de R0..R7
          ADDRin  <= 1; // habilita escrita no barramento
          DOUTin  <= 0; // não habilita escrita no barramento
          Ain     <= 0; // não carrega registrador A
          Gin     <= 0; // não carrega registrador G
          Gout    <= 0; // não lê registrador G
          Ulaop   <= 0; // não escolhe operação na ULA
          DINout  <= 0; // não coloca DIN no barramento
          Memout  <= 0; // não lê da memória
          Done    <= 0; // não indica que a instrução foi concluída
        end
      else
        begin
          // $display("[%0t] bora pic, Run = %b, Run_d = %b",$time, Run, Run_d);
          Clear   <= 0; // não limpa o contador de Tstep
          IncrPc  <= 0; // não incrementa o PC
          W_D     <= 0; // não habilita escrita na memoria
          IRin    <= 0;
          Rin     <= 8'b0;
          ADDRin  <= 0; // não habilita escrita no barramento
          DOUTin  <= 0; // não habilita escrita no barramento
          Rout    <= 8'b0;
          Ain     <= 0;
          Gin     <= 0;
          Gout    <= 0;
          Ulaop   <= 0;
          DINout  <= 0;
          Memout  <= 0; // não lê da memória
          Done    <= 0;

          case (Tstep)
            3'd0:
              begin
                // T0: carrega PC em Bus para ser escrito em Rin
                // IRin    <= 1;
                // ADDRin  <= 1; // Habilita escrita no registrador ADDR
                // Rout    <= 8'b0000_0001; // Habilita leitura do registrador PC no Bus
                // IncrPc <= 1; // Incrementa o PC se a instrução for mvi para pegar imediato
                // ADDRout
                // if (opcode == 3'b001)
                //   begin
                //   end
              end
            3'd1:
              begin
                // Rout    <= 8'b0000_0001;
                // T1: fetch da instrução na MEMORIA
                // Espera ciclo 1
              end
            3'd2:
              begin
                IRin    <= 1;
                DINout  <= 1; // Coloca DIN no barramento
                IncrPc  <= 1; // Incrementa o PC
                // ADDRin  <= 1; // Habilita escrita no barramento ADDR
              end
            3'd3:
              begin
                case (opcode)
                  mv: // mv Rx Ry
                    begin
                      Rin <= Wire_Rin; // Habilita o registrador Rx
                      Rout <= Wire_Rout; // Habilita o registrador Ry
                      Clear <= 1'b1; // Limpa o contador de Tstep
                      Done <= 1'b1; // Indica que a instrução foi concluída
                    end
                  mvi: // mvi Rx,imediato
                    begin
                      // Espera ciclo 1 para carregar o imediato da memoria
                    end
                  mvnz: // mvnz Rx,Ry
                    begin
                      Rin       <= Wire_Rin;
                      if (GRout != 0) // se G for diferente de zero
                        begin
                          Rout <= Wire_Rout; // Joga Ry em bus
                        end
                      else if (GRout == 0) // se G for igual a zero
                        begin
                          Rout <= Wire_Rin; // Joga Rx em bus (proprio dado)
                        end
                      Done      <= 1;
                      Clear     <= 1'b1; // limpa o contador de Tstep
                    end
                  add: // ADD Rx,Ry
                    begin
                      // Coloca Rout no registrador A
                      Ain  <=   1'b1;
                      Rout <=   Wire_Rin;
                    end
                  sub: // SUB Rx,Ry
                    begin
                      // Coloca Rout no registrador A
                      Ain  <=   1'b1;
                      Rout <=   Wire_Rin;
                    end
                  slt: // SLT Rx,Ry
                    begin
                      // Coloca Rout no registrador A
                      Ain  <=   1'b1;
                      Rout <=   Wire_Rin;
                    end
                  cmp: // CMP Rx,Ry
                    begin
                      // Coloca Rout no registrador A
                      Ain  <=   1'b1;
                      Rout <=   Wire_Rin;
                    end
                  ld:  // LD Rx, Ry
                    begin
                      Rout <= Wire_Rout; // Habilita o registrador Ry
                      ADDRin <= 1'b1; // Habilita escrita no barramento ADDR
                    end
                  st:  // ST Rx, Ry
                    begin
                      // Passando o dado de Rx para ser escrito na memoria
                      Rout <= Wire_Rin; // Habilita o registrador Ry
                      DOUTin <= 1'b1;   // Habilita escrita no barramento DOUT
                    end
                  push: // PUSH Rx
                    begin
                      // Fazendo $sp = $sp - 4 $sp = R6
                      Rout <= 8'b0000_0010; // Habilita o registrador R6 (SP)
                      Ulaop <= 3'b101; // Subtrai 4 na ULA
                      Gin <= 1'b1; // Habilita escrita no registrador G
                    end
                  pop: // POP Rx
                    begin
                      // Colocando SP como endereco
                      ADDRin <= 1'b1; // Habilita escrita no barramento ADDR
                      Rout <= 8'b0000_0010; // Habilita o registrador R6 (SP)
                    end
                endcase
              end
            3'd4:
              begin
                case (opcode)
                  mvi: // mvi Rx,imediato
                    begin
                      Rin <= Wire_Rin; // Habilita o registrador Rx
                      DINout <= 1'b1; // Coloca DIN no barramento
                      Done <= 1'b1; // Indica que a instrução foi concluída
                      Clear <= 1'b1; // Limpa o contador de Tstep
                      IncrPc <= 1; // Incrementa o PC pois o incremento anterior era para o imediato
                    end
                  add: // ADD Rx,Ry
                    begin
                      Rout  <= Wire_Rout; // Habilita o registrador Ry
                      Ulaop <= 3'b000;    // Subtração na ULA
                      Gin   <= 1'b1;     // Habilita escrita no registrador G
                    end
                  sub: // SUB Rx,Ry
                    begin
                      Rout  <= Wire_Rout; // Habilita o registrador Ry
                      Ulaop <= 3'b001;    // Subtração na ULA
                      Gin   <= 1'b1;     // Habilita escrita no registrador G
                    end
                  slt: // SLT Rx,Ry
                    begin
                      Rout  <= Wire_Rout; // Habilita o registrador Ry
                      Ulaop <= 3'b010;    // Set Less Than na ULA
                      Gin   <= 1'b1;     // Habilita escrita no registrador G
                    end
                  cmp: // CMP Rx,Ry
                    begin
                      Rout  <= Wire_Rout; // Habilita o registrador Ry
                      Ulaop <= 3'b011;    // Compare na ULA
                      Gin   <= 1'b1;     // Habilita escrita no registrador G
                    end
                  ld: // LD Rx,Ry
                    begin
                      // Espera 1 ciclo
                    end
                  st: // ST Rx,Ry
                    begin
                      // Passando o dado de Ry como endereco
                      Rout <= Wire_Rout; // Habilita o registrador Ry
                      ADDRin <= 1'b1; // Habilita escrita no barramento ADDR
                      W_D    <= 1'b1; // Habilita escrita no barramento DOUT
                      Done  <= 1'b1; // Indica que a instrução foi concluída
                      Clear <= 1'b1; // Limpa o contador de Tstep
                    end
                  push: // PUSH Rx
                    begin
                      // Fazendo Mem[$sp] = [Rx], $sp = R6
                      Gout   <= 1'b1; // Mandando o dado de G para o barramento
                      ADDRin <= 1'b1; // Habilita escrita no registrador ADDR 
                    end
                  pop: // POP Rx
                    begin
                      // [Rx] = Mem[$sp]
                      Rin    <= Wire_Rin; // Habilita o registrador Rx
                      Memout <= 1'b1; // Habilita leitura da memória
                    end
                endcase
              end
            3'd5:
              begin
                case (opcode)
                  add: // ADD Rx,Ry
                    begin
                      Rin   <= Wire_Rin; // Habilita o registrador Rx
                      Gout  <= 1'b1; // Habilita leitura do registrador G
                      Done  <= 1'b1; // Indica que a instrução foi concluída
                      Clear <= 1'b1; // Limpa o contador de Tstep

                      // ADD Rx,Ry
                      // Coloca Rin no bus
                      // Rout <= Wire_Rin; // Habilita o registrador Ry
                      // Gin  <= 1'b1;     // Habilita escrita no registrador G
                    end
                  sub: // SUB Rx,Ry
                    begin
                      Rin   <= Wire_Rin; // Habilita o registrador Rx
                      Gout  <= 1'b1; // Habilita leitura do registrador G
                      Done  <= 1'b1; // Indica que a instrução foi concluída
                      Clear <= 1'b1; // Limpa o contador de Tstep

                      // SUB Rx,Ry
                      // Coloca Rin no bus
                      // Rout <= Wire_Rin; // Habilita o registrador Ry
                      // Gin  <= 1'b1;     // Habilita escrita no registrador G
                    end
                  slt: // SLT Rx,Ry
                    begin
                      Rin   <= Wire_Rin; // Habilita o registrador Rx
                      Gout  <= 1'b1; // Habilita leitura do registrador G
                      Done  <= 1'b1; // Indica que a instrução foi concluída
                      Clear <= 1'b1; // Limpa o contador de Tstep
                    end
                  cmp: // CMP Rx,Ry
                    begin
                      Rin   <= Wire_Rin; // Habilita o registrador Rx
                      Gout  <= 1'b1; // Habilita leitura do registrador G
                      Done  <= 1'b1; // Indica que a instrução foi concluída
                      Clear <= 1'b1; // Limpa o contador de Tstep
                    end
                  ld: // LD Rx,Ry
                    begin
                      Rin   <= Wire_Rin; // Habilita o registrador Rx
                      Memout <= 1'b1; // Habilita leitura da memória
                      Done  <= 1'b1; // Indica que a instrução foi concluída
                      Clear <= 1'b1; // Limpa o contador de Tstep
                      // DINout <= 1'b1;    // Coloca DIN no barramento
                      // Done  <= 1'b1; // Indica que a instrução foi concluída
                      // Clear <= 1'b1; // Limpa o contador de Tstep
                      // IncrPc <= 1; // Incrementa o PC pois o incremento anterior era para o imediato
                    end
                  push: // PUSH Rx
                    begin
                      Rout   <= Wire_Rin; // Mandando o dado de Rx para o barramento
                      DOUTin <= 1'b1;     // Habilita escrita no registrador DOUT
                      W_D    <= 1'b1;     // Habilita escrita na memoria
                      Done   <= 1'b1;     // Indica que a instrução foi concluída
                      Clear  <= 1'b1;     // Limpa o contador de Tstep
                    end
                  pop: // POP Rx
                    begin
                      // Fazendo $sp = $sp + 4
                      Rout    <= 8'b0000_0010; // Escreve no registrador SP
                      Ulaop  <= 3'b100;       // Adiciona 4 na ULA
                      Gin    <= 1'b1;         // Habilita escrita no registrador G
                    end
                endcase
              end
            3'd6:
              begin
                case (opcode)
                  pop: // POP Rx
                    begin
                      // Colocando o dado de Mem[$sp] no registrador Rx
                      Rin    <= 8'b0000_0010; // Habilita escrita no registrador SP
                      Gout   <= 1'b1; // Coloca o dado de G no barramento
                      Done   <= 1'b1; // Indica que a instrução foi concluída
                      Clear  <= 1'b1; // Limpa o contador de Tstep
                    end
                endcase
              end
            // 2'b10:
            //   begin
            //     case (opcode)
            //       3'b011:
            //         begin
            //           // SUB Rx,Ry
            //           // Coloca Rin no bus
            //           Rout  <= Wire_Rout; // Habilita o registrador Ry
            //           Ulaop <= 2'b01;    // Subtração na ULA
            //           Gin   <= 1'b1;     // Habilita escrita no registrador G
            //         end
            //     endcase
            //   end

            // 2'b11:
            //   begin
            //     case (opcode)
            //       3'b011:
            //         begin
            //           Rin <= Wire_Rin; // Habilita o registrador Rx
            //           Gout <= 1'b1; // Lê o registrador G
            //           Done <= 1'b1; // Indica que a instrução foi concluída
            //           Clear <= 1'b1; // Limpa o contador de Tstep

            //           // SUB Rx,Ry
            //           // Coloca Rin no bus
            //           // Rout <= Wire_Rin; // Habilita o registrador Ry
            //           // Gin  <= 1'b1;     // Habilita escrita no registrador G
            //         end
            //     endcase
            //   end
          endcase
        end
    end


  // simples mapeamento dos campos XXX, YYY
  // supondo que você os extraia previamente em sinais separados
  // por exemplo via IR[4:6] → XXX, IR[7:9] → YYY

endmodule
