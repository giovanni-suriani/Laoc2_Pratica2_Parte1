module Pratica2_Parte1_top_level();