module unidade_controle();
  // Inputs
  input Run;
  input Resetn;

  
  // Outputs
  output Done
endmodule