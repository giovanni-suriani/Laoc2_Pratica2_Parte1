module registrador_IR(R, Rin, Clock, Q);
  // Modulo que representa um registrador de 16 bits que quando habilitado
  // armazena o valor Rin na entrada R. O valor armazenado é lido na

  // inputs
  input [8:0] R; // entrada de dados
  input Rin, Clock;

  // outputs
  output reg [8:0] Q; // valor armazenado

  // reg [8:0] Q;
  always @(posedge Clock)
    if (Rin)
      Q <= R;
endmodule
